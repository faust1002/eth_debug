module eth_debug;
endmodule
